//	logic [31:0]R2res2,R3res2;
module ForwUnitReg (R2res,R3res,R2,R3,DestR_2,DestR_3,DestR_4,R2res2,R3res2);
endmodule