module forwardMem();
endmodule