module DataMemoryTest();

	logic clk, we;
	logic[31:0] addr, wd, rd;

	DataMemory DUT(clk, we, addr, wd, rd);
	
	initial begin
		
		clk = 1'b1;
		we = 1'b0;
		addr = 32'b0;
		wd = 32'b0;
		
		#10;
		
		wd = 32'd131;
		we = 1'b1;
		clk = 1'b0;
		
		#10;
		
		clk = 1'b1;
		we = 1'b0;
		addr = 32'd1;
		wd = 32'd65;
		
		#10;
		
		clk = 1'b0;
		
		#10;
		
		addr = 32'd0;
		clk = 1'b1;
	
		#10;
	
	end

endmodule 