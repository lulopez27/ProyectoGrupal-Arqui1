module processor_tb();
	processor prcs(clk, rst);
endmodule